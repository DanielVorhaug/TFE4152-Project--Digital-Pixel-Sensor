module PIXEL_ARRAY_MEMORY_CONTROLLER (
    input logic READ_RESET,
    input logic READ_CLK,
    output logic READ_CLK_OUT,
    output logic SOMETHING_TO_POINTER //Change this name!!!
);

parameter integer WIDTH = 2;
parameter integer HEIGHT = 2;


endmodule