

module PIXEL_TOP (
    input  logic SYSTEM_CLK,
    input  logic SYSTEM_RESET,
    output logic DATA_OUT_CLK,
    output logic [OUTPUT_BUS_PIXEL_WIDTH*BIT_DEPTH-1:0] DATA_OUT
);
    
endmodule